`timescale 1ns / 1ps

module not_gate(a,b);
	input a;
	output b;
	assign b=~a;
endmodule
